`timescale 1 ps / 1 ps
module hps_driver (
        input wire                  clk,
        input wire        [7:0]     address,
        input wire                  read_en,
        output reg        [31:0]    readdata,
        input wire                  write_en,
        input wire        [31:0]    writedata,
        input wire                  chipselect,
        output reg        [7:0]     data_tx,
        output reg                  wren_fifo_tx = 1'b0,
        output reg        [7:0]     size_fifo_tx,
        input                       ready_tx,
        output reg                  start_tx = 1'b0,
        input wire        [7:0]     data_rx,
        output reg                  rden_fifo_rx = 1'b0,
        input wire        [7:0]     size_fifo_rx,
        input wire        [7:0]     interrupt_id,
        output reg                  irq = 1'b0,
        output reg                  navig_timer_start = 1'b0,
        output reg        [7:0]     led,
        output reg        [31:0]    rx_threshold = 32'd600,
        output reg        [31:0]    comp_threshold = 32'd6,
        output reg        [31:0]    guard_interval,
        output reg        [31:0]    mem_addr = 32'd0,
        input wire        [31:0]    end_address
    );

localparam  memory_size =               8'h00,
            memory_data =               8'h04,
            memory_next_tx =            8'h08,
            memory_ready =              8'h0c,
            memory_type =               8'h10,
            memory_start_tx =           8'h14,
            memory_start_navig =        8'h18,
            memory_size_rx =            8'h1c,
            memory_data_rx =            8'h20,
            memory_next_rx =            8'h24,
            memory_get_rx_threshold =   8'h28,
            memory_get_comp_threshold = 8'h2c,
            memory_get_guard_interval = 8'h30,
            memory_set_rx_threshold =   8'h34,
            memory_set_comp_threshold = 8'h38,
            memory_set_guard_interval = 8'h3c,
            memory_set_mem_addr =       8'h40,
            memory_get_end_address =    8'h44;

localparam  D_D =                   8'h01,
            N_A =                   8'h02,
            N_T =                   8'h03,
            N_Q =                   8'h04;

reg         [7:0]                   data_type = 8'd0;

always @ (posedge clk) begin

    rx_threshold <= rx_threshold ? rx_threshold : 32'd600;
    comp_threshold <= comp_threshold ? comp_threshold : 32'd6;

    if(rden_fifo_rx) begin
        rden_fifo_rx <= 1'b0;
    end
    if(wren_fifo_tx) begin
        wren_fifo_tx <= 1'b0;
    end
    if(start_tx) begin
        start_tx <= 1'b0;
    end
    if(navig_timer_start) begin
        navig_timer_start <= 1'b0;
    end
    
    if(interrupt_id) begin
        case(interrupt_id)
            D_D:
                begin
                    data_type <= D_D;
                    irq <= 1'b1;
                end

            N_A:
                begin
                    data_type <= N_A;
                    irq <= 1'b1;
                end

            N_T:
                begin
                    data_type <= N_T;
                    irq <= 1'b1;
                end

            N_Q:
                begin
                    data_tx <= N_A;
                    size_fifo_tx <= 8'd1;
                    wren_fifo_tx <= 1'b1;
                    start_tx <= 1'b1;
                end
        endcase
    end else begin
        if (chipselect) begin
            if(read_en) begin
                irq <= 1'b0;
                case(address)
                    memory_size_rx: readdata <= {24'd0, size_fifo_rx};
                    memory_data_rx: readdata <= {24'd0, data_rx};
                    memory_ready: readdata <= {31'd0, ready_tx};
                    memory_type: readdata <= {24'd0, data_type};
                    memory_get_rx_threshold: readdata <= rx_threshold;
                    memory_get_comp_threshold: readdata <= comp_threshold;
                    memory_get_guard_interval: readdata <= guard_interval;
                    memory_get_end_address: readdata <= end_address;
                endcase
            end else if(write_en) begin
                case(address)
                    memory_size: size_fifo_tx <= writedata[7:0];
                    memory_data: data_tx <= writedata[7:0];
                    memory_next_tx: wren_fifo_tx <= 1'b1;
                    memory_next_rx: rden_fifo_rx <= 1'b1;
                    memory_start_tx: start_tx <= 1'b1;
                    memory_start_navig:
                        begin
                            data_tx <= N_Q;
                            size_fifo_tx <= 8'd1;
                            wren_fifo_tx <= 1'b1;
                            navig_timer_start <= 1'b1;
                            start_tx <= 1'b1;
                        end
                    memory_set_rx_threshold: rx_threshold <= writedata;
                    memory_set_comp_threshold: comp_threshold <= writedata;
                    memory_set_guard_interval: guard_interval <= writedata;
                    memory_set_mem_addr: mem_addr <= writedata;
                endcase
            end
        end
    end
end
endmodule
