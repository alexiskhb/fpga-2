// unnamed.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module unnamed (
		output wire [12:0] streaming_source_data,  // avalon_streaming_source.data
		output wire        streaming_source_valid, //                        .valid
		input  wire        slave_clk,              //              clock_sink.clk
		input  wire        adc_clk,                //          clock_sink_adc.clk
		output wire        CONVST,                 //             conduit_end.convst
		output wire        SCK,                    //                        .sck
		output wire        SDI,                    //                        .sdi
		input  wire        SDO,                    //                        .sdo
		input  wire        slave_reset,            //              reset_sink.reset
		output wire [15:0] slave_readdata,         //                   slave.readdata
		input  wire        slave_chipselect,       //                        .chipselect
		input  wire        slave_read,             //                        .read
		input  wire        slave_address           //                        .address
	);

	adc adc_0 (
		.streaming_source_data  (streaming_source_data),  // avalon_streaming_source.data
		.streaming_source_valid (streaming_source_valid), //                        .valid
		.CONVST                 (CONVST),                 //             conduit_end.convst
		.SCK                    (SCK),                    //                        .sck
		.SDI                    (SDI),                    //                        .sdi
		.SDO                    (SDO),                    //                        .sdo
		.slave_clk              (slave_clk),              //              clock_sink.clk
		.slave_readdata         (slave_readdata),         //                   slave.readdata
		.slave_chipselect       (slave_chipselect),       //                        .chipselect
		.slave_read             (slave_read),             //                        .read
		.slave_address          (slave_address),          //                        .address
		.slave_reset            (slave_reset),            //              reset_sink.reset
		.adc_clk                (adc_clk)                 //          clock_sink_adc.clk
	);

endmodule
